module compiler_backend_vm

import rosie.parser


struct GroupBE {}

fn (mut cb GroupBE) compile(mut c Compiler, pat parser.Pattern, alias_pat parser.Pattern) ? {
	group := (alias_pat.elem as parser.GroupPattern)

	pred_p1 := c.predicate_pre(pat, 0)	// look-behind is not supported with groups

	cb.compile_inner(mut c, pat, group)?

	c.predicate_post(pat, pred_p1)
}

fn (mut cb GroupBE) compile_inner(mut c Compiler, pat parser.Pattern, group parser.GroupPattern) ? {
	add_word_boundary := group.word_boundary == true && (pat.max > 1 || pat.max == -1)

	for i in 0 .. pat.min {
		cb.compile_1(mut c, group, i > 0 && add_word_boundary)?
	}

	if pat.max != -1 {
		if pat.max > pat.min {
			for i in pat.min .. pat.max {
				cb.compile_0_or_1(mut c, group, i > 0 && add_word_boundary)?
			}
		}
	} else {
		cb.compile_0_or_many(mut c, group, add_word_boundary)?
	}
}

fn (cb GroupBE) update_addr_ar(mut c Compiler, mut ar []int, pos int) {
	for p2 in ar {
		c.update_addr(p2, c.code.len)
	}
	ar.clear()
}

fn (mut cb GroupBE) add_word_boundary(mut c Compiler) ? {
	pat := parser.Pattern{ word_boundary: false, elem: parser.NamePattern{ text: "~" }}
	c.compile_elem(pat, pat)?
}

fn (mut cb GroupBE) compile_1(mut c Compiler, group parser.GroupPattern, add_word_boundary bool) ? {
	if add_word_boundary == true { cb.add_word_boundary(mut c)? }

	mut ar := []int{}
	mut last := group.ar[0]
	for i, e in group.ar {
		if i > 0 {
			last = group.ar[i - 1]
			if last.operator == .choice  {
				// Wrap every choice ...
				p1 := c.add_choice(0)
				c.compile_elem(e, e)?
				ar << c.add_commit(0)	// pop the entry added by choice	// TODO Not sure commit is the right thin to do here
				c.update_addr(p1, c.code.len)
			} else if last.operator == .sequence {
				// End of choices
				if ar.len > 0 {
					c.add_fail()
					cb.update_addr_ar(mut c, mut ar, c.code.len)
				}

				if last.word_boundary == true { cb.add_word_boundary(mut c)? }
				c.compile_elem(e, e)?
			} else {
				panic("GroupBE: compile_1: unsupported construct: ${group.repr()}")
			}
		} else if e.operator == .choice {
			// Wrap every choice ...
			p1 := c.add_choice(0)
			c.compile_elem(e, e)?
			ar << c.add_commit(0)	// pop the entry added by choice	// TODO Not sure commit is the right thin to do here
			c.update_addr(p1, c.code.len)
		} else if e.operator == .sequence {
			c.compile_elem(e, e)?
		} else {
			panic("GroupBE: compile_1: unsupported construct: ${group.repr()}")
		}
	}

	if ar.len > 0 {
		c.add_fail()
		cb.update_addr_ar(mut c, mut ar, c.code.len)
	}
}

fn (mut cb GroupBE) compile_0_or_many(mut c Compiler, group parser.GroupPattern, add_word_boundary bool) ? {
	p1 := c.add_choice(0)
	p2 := c.code.len
	cb.compile_1(mut c, group, add_word_boundary)?
	c.add_partial_commit(p2)
	c.update_addr(p1, c.code.len)
}

fn (mut cb GroupBE) compile_1_or_many(mut c Compiler, group parser.GroupPattern, add_word_boundary bool) ? {
	cb.compile_1(mut c, group, add_word_boundary)?
	cb.compile_0_or_many(mut c, group, add_word_boundary)?
}

fn (mut cb GroupBE) compile_0_or_1(mut c Compiler, group parser.GroupPattern, add_word_boundary bool) ? {
	p1 := c.add_choice(0)
	cb.compile_1(mut c, group, add_word_boundary)?
	p2 := c.add_commit(0)	// TODO Not sure commit is the right thin to do here
	c.update_addr(p1, c.code.len)
	c.update_addr(p2, c.code.len)
}
