module vlang

// This file is copied 1:1 to the generate module

fn test_dummy() ? {
	// Only to test successful compilation
	assert true
}