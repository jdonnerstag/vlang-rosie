module stage_0

// This is the module description for parser_stage_0. A handwritten parser to bootstrap
// vrosie.
