module compiler_backend_vm

import rosie.parser


struct DisjunctionBE {
pub:
	pat parser.Pattern
	elem parser.DisjunctionPattern
}


fn (cb DisjunctionBE) compile(mut c Compiler) ? {
	mut x := DefaultPatternCompiler{
		pat: cb.pat,
		predicate_be: DefaultPredicateBE{ pat: cb.pat },
		compile_1_be: cb,
		compile_0_to_many_be: DefaultCompile_0_to_many{ pat: cb.pat, compile_1_be: cb }
	}

	x.compile(mut c) ?
}

fn (cb DisjunctionBE) compile_1(mut c Compiler) ? {
	group := cb.elem
	if group.negative == false {
		mut ar := []int{}
		for i, e in group.ar {
			if (i + 1) == group.ar.len {
				c.compile_elem(e, e)?
			} else {
				// Some pattern can be performance optimized by avoiding .choice
				// TODO Identify additional pattern that may benefit from it. Charsets?
				if e.elem is parser.LiteralPattern {
					str := e.elem.text
					if str.len > 0 {
						p2 := c.add_test_char(str[0], 0)
						mut ee := e
						ee.elem = parser.LiteralPattern{ text: str[1 ..] }
						p1 := c.add_choice(0)
						c.add_any()
						c.compile_elem(ee, ee)?
						ar << c.add_commit(0)
						c.update_addr(p1, c.code.len)
						c.update_addr(p2, c.code.len)
					}
				} else {
					p1 := c.add_choice(0)
					c.compile_elem(e, e)?
					ar << c.add_commit(0)
					c.update_addr(p1, c.code.len)
				}
			}
		}

		for p2 in ar { c.update_addr(p2, c.code.len) }
	} else {
		for e in group.ar {
			p1 := c.add_choice(0)
			c.compile_elem(e, e)?
			p2 := c.add_commit(0)
			p3 := c.add_fail()
			c.update_addr(p2, p3)
			c.update_addr(p1, c.code.len)
		}

		c.add_any()
	}
}
