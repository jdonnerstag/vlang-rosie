module mytest

fn test_dummy() ? {
	// Only to test successful compilation
	assert true
}