module rpl_3_0

fn test_import() ? {
	// RPL 3.0 does not support the grammar syntax any longer
}

fn test_grammar_stmt() ? {
	// RPL 3.0 does not support the grammar syntax any longer
}
/* */