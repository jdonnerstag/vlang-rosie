module rpl

import os


fn (mut p Parser) find_rpl_file(name string) ? string {
	if name.ends_with(".rpl") {
		return p.find_rpl_file(name[0 .. name.len - 4])
	}

	if name.len == 0 {
		return error("Import name must not be empty. File=$name")
	}

	for path in p.import_path {
		if f := p.find_rpl_file_("${path}/${name}") {
			return f
		}
	}

	if f := p.find_rpl_file_(name) {
		return f
	}

	return error("Import package: File not found: name='$name', path=${p.import_path}. ")
}

fn (mut p Parser) find_rpl_file_(name string) ? string {
	if os.is_file(name) {
		return os.real_path(name)
	}

	fp := "${name}.rpl"
	if os.is_file(fp) {
		return os.real_path(fp)
	}

	return none
}

fn (mut p Parser) find_and_load_package(name string) ?string {
	fpath := p.find_rpl_file(name)?
	eprintln("fpath: $fpath")

	if p.package_cache.contains(fpath) {
		eprintln("Package has already been imported: $fpath")
		return fpath
	}

	if p.debug > 10 {
		eprintln(">> Import: load and parse '$fpath'")
		defer { eprintln("<< Import: load and parse '$fpath'") }
	}

	mut p2 := p.clone()
	p2.parse(file: fpath) or {
		return error("${err.msg}; file: $fpath")
	}

	p2.main.name = if p2.package.len > 0 { p2.package } else { name }
	p2.main.fpath = fpath
	eprintln("Add package to cache: $p2.main.name, $p2.main.fpath")
	p2.package_cache.add_package(p2.main)?	// TODO may be rename add_package() to add(). Though add_package() can be found more easily

	return fpath
}

fn (mut p Parser) import_package(alias string, name string) ? {
	eprintln("import_package: '$name'")
	fpath := p.find_and_load_package(name) or {
		return error("RPL parser: Failed to import package '$name': $err.msg")
	}
	eprintln("Import package: alias: '$alias', name: '$name', fpath: '$fpath'")
	p.package().imports[alias] = fpath
}
