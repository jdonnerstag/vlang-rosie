
module rosie

pub struct Engine {
pub:
	debug int

pub mut:
	package_cache 	 PackageCache
//	parser 			 parser.Parser
	// optimizer OptimizerInterface
	// compiler CompilerInterface
	// runtime RuntimeInterface
}
