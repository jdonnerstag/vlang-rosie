module v2

// The only purpose for this file is to make sure that the V2 runtime
// compiles successfully.

fn test_simple_00() ? {
}
/* */