module vm_v2

import rosie
import rosie.runtimes.v2 as rt

struct Compiler {
pub:
	unit_test bool				// When compiling for unit tests, then capture ALL variables (incl. alias)

pub mut:
	current &rosie.Package		// The current package context: either "main" or a grammar package
	rplx &rosie.Rplx				// symbols, charsets, instructions
	func_implementations map[string]int		// function name => pc: fn entry point
	debug int
	indent_level int
	user_captures []string		// User may override which variables are captured. (back-refs are always captured)
}

[params]
pub struct FnNewCompilerOptions {
pub:
	rplx &rosie.Rplx = rosie.new_rplx()
	user_captures []string
	unit_test bool
	debug int
	indent_level int = 2
}

pub fn new_compiler(main &rosie.Package, args FnNewCompilerOptions) ? Compiler {
	return Compiler{
		current: main
		rplx: args.rplx
		debug: args.debug
		indent_level: args.indent_level
		unit_test: args.unit_test
		user_captures: args.user_captures
	}
}

pub fn (c Compiler) input_len(pat rosie.Pattern) ? int {
	if pat.elem is rosie.NamePattern {
		b := c.current.get(pat.elem.name)?
		if b.grammar.len > 0 {
			return none	  // Unable to determine input length for recursive pattern
		}
		return c.input_len(b.pattern)
	} else if pat.elem is rosie.GroupPattern {
		// TODO: GroupPattern has an input_len() method, but it is not able to resolve NamePattern.
		mut len := 0
		for p in pat.elem.ar {
			if p.predicate != .na {
				len += c.input_len(p) or {
					return err
				}
			}
		}
		return len
	}

	// Ignore the predicate of the outer most pattern, because it is the input-len
	// of this pattern, that we want to determine.
	return pat.elem.input_len()
}

// compile Compile the necessary instructions for a specific
// (public) binding from the rpl file. Use "*" for anonymous
// pattern.
pub fn (mut c Compiler) compile(name string) ? {
	// Set the context used to resolve variable names
	orig_current := c.current
	defer { c.current = orig_current }

	if c.debug > 0 { eprintln("Compile pattern for binding='$name'") }
	b, new_current := c.current.get_bp(name)?
	c.current = new_current
	if c.debug > 0 { eprintln("Compile: current='${new_current.name}'; ${b.repr()}") }

	//eprintln("Compiler: name='$name', package='$b.package', grammar='$b.grammar', current='$c.current.name', repr=${b.pattern.repr()}")
	// ------------------------------------------

	if b.recursive == true || b.func == true {
		c.compile_func_body(b)?
	}

	full_name := b.full_name()
	c.rplx.entrypoints.add(name: full_name, start_pc: c.rplx.code.len)?

	pat := b.pattern
	if func_pc := c.func_implementations[full_name] {
		c.add_call(func_pc, full_name)
	} else {
		c.add_open_capture(full_name)
		c.compile_elem(pat, pat)?
		c.add_close_capture()
	}
	c.add_end()
}

pub fn (mut c Compiler) compile_func_body(b rosie.Binding) ? {
	full_name := b.full_name()
	if full_name in c.func_implementations {
		return
	}

	if b.recursive { c.add_register_recursive(full_name) }

	mut p1 := c.add_jmp(0)
	c.func_implementations[full_name] = c.rplx.code.len

	add_capture := b.alias == false || c.unit_test
	if add_capture { c.add_open_capture(full_name) }

	p2 := c.add_choice(0)

	c.compile_elem(b.pattern, b.pattern)?

	if add_capture { c.add_close_capture() }

	c.add_ret()
	c.update_addr(p2, c.rplx.code.len)
	c.add_fail_twice()
	c.update_addr(p1, c.rplx.code.len)
}

fn (mut c Compiler) compile_elem(pat rosie.Pattern, alias_pat rosie.Pattern) ? {
	//eprintln("compile_elem: ${pat.repr()}")
	mut be := PatternCompiler(StringBE{})

	match pat.elem {
		rosie.LiteralPattern { be = PatternCompiler(StringBE{ pat: pat, text: pat.elem.text }) }
		rosie.CharsetPattern { be = PatternCompiler(CharsetBE{ pat: pat, cs: pat.elem.cs }) }
		rosie.GroupPattern { be = PatternCompiler(GroupBE{ pat: pat, elem: pat.elem }) }
		rosie.DisjunctionPattern { be = PatternCompiler(DisjunctionBE{ pat: pat, elem: pat.elem }) }
		rosie.NamePattern { be = PatternCompiler(AliasBE{ pat: pat, name: pat.elem.name }) }
		rosie.EofPattern { be = PatternCompiler(EofBE{ pat: pat, eof: pat.elem.eof }) }
		rosie.MacroPattern { be = PatternCompiler(MacroBE{ pat: pat, elem: pat.elem }) }
		rosie.FindPattern { be = PatternCompiler(FindBE{ pat: pat, elem: pat.elem }) }
		rosie.NonePattern { return error("Pattern not initialized !!!") }
	}

	be.compile(mut c)?
}

pub fn (mut c Compiler) add_open_capture(name string) int {
	idx := c.rplx.symbols.add(name)
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.open_capture).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_behind(offset int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.behind).set_aux(offset))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_close_capture() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.close_capture))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_end() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.end))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_digit() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.digit))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_ret() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.ret))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_fail() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.fail))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_fail_twice() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.fail_twice))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_test_any(pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.test_any))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_char(ch byte) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.char).set_char(ch))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_until_char(ch byte, fail bool) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.until_char).set_char(ch))
	c.rplx.code << rosie.Slot(if fail { u32(0) } else { u32(-1) })
	return rtn
}

pub fn (mut c Compiler) add_span(cs rosie.Charset) int {
	idx := c.rplx.add_cs(cs)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.span).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_test_char(ch byte, pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.test_char).set_char(ch))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_if_char(ch byte, pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.if_char).set_char(ch))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_choice(pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.choice))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_partial_commit(pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.partial_commit))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_back_commit(pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.back_commit))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_any() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.any))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_commit(pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.commit))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_call(fn_pos int, fn_name string) int {
	idx := c.rplx.symbols.add(fn_name)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.call).set_aux(idx))
	c.rplx.code << fn_pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_jmp(pos int) int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.jmp))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_set(cs rosie.Charset) int {
	idx := c.rplx.add_cs(cs)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.set).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_until_set(cs rosie.Charset, fail bool) int {
	idx := c.rplx.add_cs(cs)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.until_set).set_aux(idx))
	c.rplx.code << rosie.Slot(if fail { u32(0) } else { u32(-1) })
	return rtn
}

pub fn (mut c Compiler) add_test_set(cs rosie.Charset, pos int) int {
	idx := c.rplx.add_cs(cs)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.test_set).set_aux(idx))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_if_str(str string, pos int) int {
	idx := c.rplx.symbols.add(str)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.if_str).set_aux(idx))
	c.rplx.code << pos - rtn
	return rtn
}

pub fn (mut c Compiler) add_str(str string) int {
	idx := c.rplx.symbols.add(str)

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.str).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_message(str string) int {
	idx := c.rplx.symbols.add(str)
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.message).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_backref(name string) ? int {
	idx := c.rplx.symbols.find(name) or {
		return error("Unable to find back-referenced binding in symbol table: '$name'")
	}

	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.backref).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_register_recursive(name string) int {
	idx := c.rplx.symbols.add(name)
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.register_recursive).set_aux(idx))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_word_boundary() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.word_boundary))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_dot_instr() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.dot))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_bit_7() int {
	rtn := c.rplx.code.len
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.bit_7))
	c.rplx.code << rosie.Slot(0)
	return rtn
}

pub fn (mut c Compiler) add_quote(ch1 byte, ch2 byte, esc byte, stop byte) int {
	rtn := c.rplx.code.len
	mut data := u32(0)
	unsafe {
		mut ptr := &byte(&data)
		ptr[0] = ch1
		ptr[1] = ch2
		ptr[2] = esc
		ptr[3] = stop
	}
	c.rplx.code << rosie.Slot(rt.opcode_to_bytecode(.quote))
	c.rplx.code << rosie.Slot(data)
	return rtn
}

pub fn (mut c Compiler) update_addr(pc int, pos int) {
	c.rplx.code[pc + 1] = pos - pc
}
