module rpl_1_3

// This is the module description for parser_rpl. A parser that uses vrosie to parse
// rpl-files and rpl-pattern. This is the default parser under normal circumstances.
