// ----------------------------------------------------------------------------
// Analyze the AST of a single pattern and optimize it
// ----------------------------------------------------------------------------

module parser

fn (mut parser Parser) optimize(pattern Pattern) Pattern {
	return pattern
}
