module rpl_3_0

// A RPL-3.0 parser, leveraging RPL-1.3 to create the parser.