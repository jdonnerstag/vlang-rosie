module core_0

// This is the module description for parser_core_0. A handwritten parser to bootstrap
// vrosie.
